		
	

	



