module clkrst (clk, rst_n);

    output reg clk;
    output reg rst_n;

    initial begin

	  

	  
    end



endmodule
