module uart_TX(
    input	      clk,                  //系统时钟
    input         rst_n,                //系统复位，低电平有效
    
    input         uart_en,                  //发送使能信号
    input  [7:0]  uart_din,                 //待发送数据
    output  reg   TX,                  //UART发送端口
	output		  tx_done
    );
    
//parameter define
parameter  CLK_FREQ = 50000000;             //系统时钟频率
parameter  UART_BPS = 115200;                 //串口波特率
localparam BPS_CNT  = CLK_FREQ/UART_BPS;    //为得到指定波特率，对系统时钟计数BPS_CNT次

//reg define
reg        uart_en_d0; 
reg        uart_en_d1;  
reg [15:0] clk_cnt;                         //系统时钟计数器
reg [ 3:0] tx_cnt;                          //发送数据计数器
reg        tx_flag;                         //发送过程标志信号
reg [ 7:0] tx_data;                         //寄存发送数据

//wire define
wire       en_flag;

//*****************************************************
//**                    main code
//*****************************************************
//捕获uart_en上升沿，得到一个时钟周期的脉冲信号
assign en_flag = (~uart_en_d1) & uart_en_d0;

//negedge for tx_flag means tx done
reg dff1, dff2;
always @ (posedge clk, negedge rst_n) begin
	if (!rst_n) begin
		dff1 <= 1'b0;
		dff2 <= 1'b0;
	end else begin
		dff1 <= tx_flag;
		dff2 <= dff1;
	end
end
assign tx_done = (!dff1) & (dff2);
                                                 
//对发送使能信号uart_en延迟两个时钟周期
always @(posedge clk or negedge rst_n) begin         
    if (!rst_n) begin
        uart_en_d0 <= 1'b0;                                  
        uart_en_d1 <= 1'b0;
    end                                                      
    else begin                                               
        uart_en_d0 <= uart_en;                               
        uart_en_d1 <= uart_en_d0;                            
    end
end

//当脉冲信号en_flag到达时,寄存待发送的数据，并进入发送过程          
always @(posedge clk or negedge rst_n) begin         
    if (!rst_n) begin                                  
        tx_flag <= 1'b0;
        tx_data <= 8'd0;
    end 
    else if (en_flag) begin                 //检测到发送使能上升沿                      
            tx_flag <= 1'b1;                //进入发送过程，标志位tx_flag拉高
            tx_data <= uart_din;            //寄存待发送的数据
        end
        else 
        //if ((tx_cnt == 4'd9)&&(clk_cnt == BPS_CNT/2))
		if ((tx_cnt == 4'd9)&&(clk_cnt == BPS_CNT-1))
        begin                               //计数到停止位中间时，停止发送过程
            tx_flag <= 1'b0;                //发送过程结束，标志位tx_flag拉低
            tx_data <= 8'd0;
        end
        else begin
            tx_flag <= tx_flag;
            tx_data <= tx_data;
        end 
end

//进入发送过程后，启动系统时钟计数器与发送数据计数器
always @(posedge clk or negedge rst_n) begin         
    if (!rst_n) begin                             
        clk_cnt <= 16'd0;                                  
        tx_cnt  <= 4'd0;
    end                                                      
    else if (tx_flag) begin                 //处于发送过程
        if (clk_cnt < BPS_CNT - 1) begin
            clk_cnt <= clk_cnt + 1'b1;
            tx_cnt  <= tx_cnt;
        end
        else begin
            clk_cnt <= 16'd0;               //对系统时钟计数达一个波特率周期后清零
            tx_cnt  <= tx_cnt + 1'b1;       //此时发送数据计数器加1
        end
    end
    else begin                              //发送过程结束
        clk_cnt <= 16'd0;
        tx_cnt  <= 4'd0;
    end
end

//根据发送数据计数器来给uart发送端口赋值
always @(posedge clk or negedge rst_n) begin        
    if (!rst_n)  
        TX <= 1'b1;        
    else if (tx_flag)
        case(tx_cnt)
            4'd0: TX <= 1'b0;         //起始位 
            4'd1: TX <= tx_data[0];   //数据位最低位
            4'd2: TX <= tx_data[1];
            4'd3: TX <= tx_data[2];
            4'd4: TX <= tx_data[3];
            4'd5: TX <= tx_data[4];
            4'd6: TX <= tx_data[5];
            4'd7: TX <= tx_data[6];
            4'd8: TX <= tx_data[7];   //数据位最高位
            4'd9: TX <= 1'b1;         //停止位
            default: ;
        endcase
    else 
        TX <= 1'b1;                   //空闲时发送端口为高电平
end

endmodule	          