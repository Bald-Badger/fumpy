`include "../param.vh"

module systolic_arr_ctrl (
	
);

endmodule
